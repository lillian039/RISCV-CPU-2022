module branch_target_buffer('
);
endmodule
